--
-- VHDL Architecture my_project4_lib.merge.rtl
--
-- Created:
--          by - ELHUSSEIN-STORE.UNKNOWN (DESKTOP-NC58NV1)
--          at - 17:20:22 04/28/2025
--
-- using Mentor Graphics HDL Designer(TM) 2021.1 Built on 14 Jan 2021 at 15:11:42
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY merge IS
  port(a,b: in std_logic_vector(3 downto 0);
  z:out std_logic_vector(7 downto 0));
END ENTITY merge;

--
ARCHITECTURE rtl OF merge IS
BEGIN
  z<= a&b;
END ARCHITECTURE rtl;

