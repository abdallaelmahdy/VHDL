--
-- VHDL Architecture my_project4_lib.and_4.rtl
--
-- Created:
--          by - ELHUSSEIN-STORE.UNKNOWN (DESKTOP-NC58NV1)
--          at - 04:15:13 04/28/2025
--
-- using Mentor Graphics HDL Designer(TM) 2021.1 Built on 14 Jan 2021 at 15:11:42
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY and_4 IS
  port(a,b: in std_logic;
  y:out std_logic);
END ENTITY and_4;

--
ARCHITECTURE rtl OF and_4 IS
BEGIN
  y<= (a AND b);
END ARCHITECTURE rtl;

